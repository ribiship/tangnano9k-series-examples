module oled(
    input clk,
    input btn1,
    input btn2,
    output [5:0] led
);
